library verilog;
use verilog.vl_types.all;
entity MAC_to_maddr_tb is
end MAC_to_maddr_tb;
