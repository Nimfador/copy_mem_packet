// Vozmozhno, sdelat' bufer kol'tsevim
module reg_file
    #(
        parameter               pBITS = 8,      //Data Width
                                pWIDHT = 3072   //Number of regs or depth of data
    )
    (
        input wire              iclk,
        input wire              iwr_en,
        input wire [pWIDHT-1:0] iw_addr,
        input wire [pWIDHT-1:0] ir_addr,
        input wire [pBITS-1:0]  iw_reg_data,
        output wire [pBITS-1:0] or_data
    );

    // signal declaration
    reg [pBITS-1:0] rarray [pWIDHT-1:0];
    
    // body
    always @(posedge iclk ) begin
        if (iwr_en) begin                           // write
            rarray[iw_addr] <= iw_reg_data;    
        end
      
    end

    assign or_data = rarray[ir_addr];

endmodule