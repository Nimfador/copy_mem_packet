module FSM_mem_read 
    #(
        parameter pPORT_NUM = 4,
    )(
        input wire [$clog2(pPORT_NUM)-1:0]
    );

endmodule
