library verilog;
use verilog.vl_types.all;
entity Ethernet_RX_frame_analyzer_tb is
end Ethernet_RX_frame_analyzer_tb;
