library verilog;
use verilog.vl_types.all;
entity crc_v_unit is
end crc_v_unit;
