library verilog;
use verilog.vl_types.all;
entity project_header_v_unit is
end project_header_v_unit;
