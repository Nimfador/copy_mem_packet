library verilog;
use verilog.vl_types.all;
entity copy_packet_to_mem_tb is
end copy_packet_to_mem_tb;
