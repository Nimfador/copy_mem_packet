library verilog;
use verilog.vl_types.all;
entity FSM_frame_vlg_tst is
end FSM_frame_vlg_tst;
