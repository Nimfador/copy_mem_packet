library verilog;
use verilog.vl_types.all;
entity copy_packet_to_mem_sv_unit is
end copy_packet_to_mem_sv_unit;
